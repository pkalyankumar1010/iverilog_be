module test; 
initial begin 
$display("Hello, Verilog");
end endmodule