module test; 
initial begin
$display("Hello, 3 Verilog");
end endmodule